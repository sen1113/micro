module flags();

endmodule
