module mdr();

endmodule
