module dr();

endmodule
