`define f 4
`define r 3
`define x 2
`define m 1
`define w 0

module  register_file(ra1, ra2, wa, rd1, rd2, wd, we, clk, n_rst//, rf
);
	input  [ 2:0] ra1, ra2, wa;	// �A�h���X�i���W�X�^�ԍ��j
	output [31:0] rd1, rd2;    	// �ǂݏo���f�[�^
	input  [31:0] wd;         	// �������݃f�[�^
	input  we;                  	// ���C�g�E�C�l�[�u��
	input  clk, n_rst;         	// �N���b�N�C���Z�b�g
     // output reg [31:0] rf[0:7];	// ���W�X�^�E�t�@�C���{�́i�f�o�O�p�o�́j

 	integer i;

	reg [31:0] rf [0:7];        	// 32-bit x 8-word ���W�X�^�E�t�@�C���{��
	always @(posedge clk  or  negedge n_rst) begin
	   if (n_rst == 0)
	        for (i = 0; i < 8; i = i + 1)
	            rf[i] <= 0;
	   else if (we == 1) 
	        rf[wa] <= wd;        	// ��������
	end

	assign  rd1 = rf[ra1];  	// �ǂݏo��
	assign  rd2 = rf[ra2];  	// �ǂݏo��

endmodule