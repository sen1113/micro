module alu();

endmodule
